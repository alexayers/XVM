/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
MATH.VH
Math Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/

function float cos(float flt);

function float sin(float flt);

function float tan(float flt);

function float acos(float flt);

function float asin(float flt);

function float atan(float flt);

function float atan2(float x, float y);

function float cosh(float flt);

function float sinh(float flt);

function float tanh(float flt);

function float exp(float flt);

function float log(float flt);

function float log10(float flt);

function float pow(float base,float exponent);

function float sqrt(float flt);

function float ceil(float flt);

function float fabs(float flt);

function float floor(float flt);