/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
STRING.VH
String Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/

function int strlen(string str);
//Returns lenght of string.

function string substr(string str, int start, int end);
//Returns a substring

function string strtolower(string str);
//Returns all lowercase string.

function string strtoupper(string str);
//Returns all uppercase string.

function string strreplace(string str, string find, string replace);
//Replaces substring within a string with another string.

function int strstr(string str, string haystack, string needle);








