/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
DEBUG.VH
Debug Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/

 