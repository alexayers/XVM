/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
SOCKET.VH
Networking Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/






