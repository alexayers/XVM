/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
SYSTEM.VH
System Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/

function int tickcount();
//Returns native system tickcount.

function string osinfo();
//Returns operation system information.

function string meminfo();
//Returns memory information.

function string cpuinfo();
//Returns cpu information.




