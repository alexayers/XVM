/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
DATE.VH
Date & Time Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/

function string time();

function string date();

function int hour();

function int minute();

function int second();

function int millisecond();

function int ampm();

function int month();

function int day();

function int year();

