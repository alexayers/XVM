/*
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
STDLIB.VH
Standard Library
Developed by: Alex Ayers
AYERSLABS 2009
-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-=-
*/

function int atoi(string str);
//ASCII to Integer

function string itoa(int num);
//Integer to ASCII

function string ftoa(float num);
//Float to ASCII

function float itof(int num);
//Integer to Float

function float stof(int num);
//String to Float

function int rand();
//Generates a random number.

function void sleep(int milliseconds);
//Pauses program execution for specified number of milliseconds.

function void exit();
